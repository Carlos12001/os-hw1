// cpu.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module cpu (
		input  wire       clk_clk,                                    //                                 clk.clk
		output wire [7:0] leds_minutes_ls_external_connection_export, // leds_minutes_ls_external_connection.export
		output wire [7:0] leds_minutes_ms_external_connection_export, // leds_minutes_ms_external_connection.export
		output wire [6:0] leds_seconds_ls_external_connection_export, // leds_seconds_ls_external_connection.export
		output wire [6:0] leds_seconds_ms_external_connection_export, // leds_seconds_ms_external_connection.export
		input  wire       pio_key_0_external_connection_export,       //       pio_key_0_external_connection.export
		input  wire       pio_key_1_external_connection_export,       //       pio_key_1_external_connection.export
		input  wire       pio_key_2_external_connection_export,       //       pio_key_2_external_connection.export
		input  wire       pio_key_3_external_connection_export,       //       pio_key_3_external_connection.export
		input  wire [1:0] pio_switches_external_connection_export,    //    pio_switches_external_connection.export
		input  wire       reset_reset_n                               //                               reset.reset_n
	);

	wire  [31:0] cpu_data_master_readdata;                                    // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                 // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                 // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [19:0] cpu_data_master_address;                                     // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                  // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                        // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                       // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                   // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                             // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                          // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [19:0] cpu_instruction_master_address;                              // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                 // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;              // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;           // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;           // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;               // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                  // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;            // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                 // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;             // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_memoria_s1_chipselect;                     // mm_interconnect_0:memoria_s1_chipselect -> memoria:chipselect
	wire  [31:0] mm_interconnect_0_memoria_s1_readdata;                       // memoria:readdata -> mm_interconnect_0:memoria_s1_readdata
	wire   [9:0] mm_interconnect_0_memoria_s1_address;                        // mm_interconnect_0:memoria_s1_address -> memoria:address
	wire   [3:0] mm_interconnect_0_memoria_s1_byteenable;                     // mm_interconnect_0:memoria_s1_byteenable -> memoria:byteenable
	wire         mm_interconnect_0_memoria_s1_write;                          // mm_interconnect_0:memoria_s1_write -> memoria:write
	wire  [31:0] mm_interconnect_0_memoria_s1_writedata;                      // mm_interconnect_0:memoria_s1_writedata -> memoria:writedata
	wire         mm_interconnect_0_memoria_s1_clken;                          // mm_interconnect_0:memoria_s1_clken -> memoria:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                       // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                         // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                          // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                            // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                        // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_leds_seconds_ls_s1_chipselect;             // mm_interconnect_0:leds_seconds_ls_s1_chipselect -> leds_seconds_ls:chipselect
	wire  [31:0] mm_interconnect_0_leds_seconds_ls_s1_readdata;               // leds_seconds_ls:readdata -> mm_interconnect_0:leds_seconds_ls_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_seconds_ls_s1_address;                // mm_interconnect_0:leds_seconds_ls_s1_address -> leds_seconds_ls:address
	wire         mm_interconnect_0_leds_seconds_ls_s1_write;                  // mm_interconnect_0:leds_seconds_ls_s1_write -> leds_seconds_ls:write_n
	wire  [31:0] mm_interconnect_0_leds_seconds_ls_s1_writedata;              // mm_interconnect_0:leds_seconds_ls_s1_writedata -> leds_seconds_ls:writedata
	wire         mm_interconnect_0_leds_seconds_ms_s1_chipselect;             // mm_interconnect_0:leds_seconds_ms_s1_chipselect -> leds_seconds_ms:chipselect
	wire  [31:0] mm_interconnect_0_leds_seconds_ms_s1_readdata;               // leds_seconds_ms:readdata -> mm_interconnect_0:leds_seconds_ms_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_seconds_ms_s1_address;                // mm_interconnect_0:leds_seconds_ms_s1_address -> leds_seconds_ms:address
	wire         mm_interconnect_0_leds_seconds_ms_s1_write;                  // mm_interconnect_0:leds_seconds_ms_s1_write -> leds_seconds_ms:write_n
	wire  [31:0] mm_interconnect_0_leds_seconds_ms_s1_writedata;              // mm_interconnect_0:leds_seconds_ms_s1_writedata -> leds_seconds_ms:writedata
	wire         mm_interconnect_0_leds_minutes_ls_s1_chipselect;             // mm_interconnect_0:leds_minutes_ls_s1_chipselect -> leds_minutes_ls:chipselect
	wire  [31:0] mm_interconnect_0_leds_minutes_ls_s1_readdata;               // leds_minutes_ls:readdata -> mm_interconnect_0:leds_minutes_ls_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_minutes_ls_s1_address;                // mm_interconnect_0:leds_minutes_ls_s1_address -> leds_minutes_ls:address
	wire         mm_interconnect_0_leds_minutes_ls_s1_write;                  // mm_interconnect_0:leds_minutes_ls_s1_write -> leds_minutes_ls:write_n
	wire  [31:0] mm_interconnect_0_leds_minutes_ls_s1_writedata;              // mm_interconnect_0:leds_minutes_ls_s1_writedata -> leds_minutes_ls:writedata
	wire         mm_interconnect_0_leds_minutes_ms_s1_chipselect;             // mm_interconnect_0:leds_minutes_ms_s1_chipselect -> leds_minutes_ms:chipselect
	wire  [31:0] mm_interconnect_0_leds_minutes_ms_s1_readdata;               // leds_minutes_ms:readdata -> mm_interconnect_0:leds_minutes_ms_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_minutes_ms_s1_address;                // mm_interconnect_0:leds_minutes_ms_s1_address -> leds_minutes_ms:address
	wire         mm_interconnect_0_leds_minutes_ms_s1_write;                  // mm_interconnect_0:leds_minutes_ms_s1_write -> leds_minutes_ms:write_n
	wire  [31:0] mm_interconnect_0_leds_minutes_ms_s1_writedata;              // mm_interconnect_0:leds_minutes_ms_s1_writedata -> leds_minutes_ms:writedata
	wire  [31:0] mm_interconnect_0_pio_switches_s1_readdata;                  // pio_switches:readdata -> mm_interconnect_0:pio_switches_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_switches_s1_address;                   // mm_interconnect_0:pio_switches_s1_address -> pio_switches:address
	wire  [31:0] mm_interconnect_0_pio_key_0_s1_readdata;                     // pio_key_0:readdata -> mm_interconnect_0:pio_key_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_key_0_s1_address;                      // mm_interconnect_0:pio_key_0_s1_address -> pio_key_0:address
	wire  [31:0] mm_interconnect_0_pio_key_1_s1_readdata;                     // pio_key_1:readdata -> mm_interconnect_0:pio_key_1_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_key_1_s1_address;                      // mm_interconnect_0:pio_key_1_s1_address -> pio_key_1:address
	wire  [31:0] mm_interconnect_0_pio_key_2_s1_readdata;                     // pio_key_2:readdata -> mm_interconnect_0:pio_key_2_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_key_2_s1_address;                      // mm_interconnect_0:pio_key_2_s1_address -> pio_key_2:address
	wire         mm_interconnect_0_pio_key_3_s1_chipselect;                   // mm_interconnect_0:pio_key_3_s1_chipselect -> pio_key_3:chipselect
	wire  [31:0] mm_interconnect_0_pio_key_3_s1_readdata;                     // pio_key_3:readdata -> mm_interconnect_0:pio_key_3_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_key_3_s1_address;                      // mm_interconnect_0:pio_key_3_s1_address -> pio_key_3:address
	wire         mm_interconnect_0_pio_key_3_s1_write;                        // mm_interconnect_0:pio_key_3_s1_write -> pio_key_3:write_n
	wire  [31:0] mm_interconnect_0_pio_key_3_s1_writedata;                    // mm_interconnect_0:pio_key_3_s1_writedata -> pio_key_3:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // pio_key_3:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_irq_irq;                                                 // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [cpu:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, leds_minutes_ls:reset_n, leds_minutes_ms:reset_n, leds_seconds_ls:reset_n, leds_seconds_ms:reset_n, memoria:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, pio_key_0:reset_n, pio_key_1:reset_n, pio_key_2:reset_n, pio_key_3:reset_n, pio_switches:reset_n, rst_translator:in_reset, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [cpu:reset_req, memoria:reset_req, rst_translator:reset_req_in]

	cpu_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	cpu_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	cpu_leds_minutes_ls leds_minutes_ls (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_leds_minutes_ls_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_minutes_ls_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_minutes_ls_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_minutes_ls_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_minutes_ls_s1_readdata),   //                    .readdata
		.out_port   (leds_minutes_ls_external_connection_export)       // external_connection.export
	);

	cpu_leds_minutes_ls leds_minutes_ms (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_leds_minutes_ms_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_minutes_ms_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_minutes_ms_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_minutes_ms_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_minutes_ms_s1_readdata),   //                    .readdata
		.out_port   (leds_minutes_ms_external_connection_export)       // external_connection.export
	);

	cpu_leds_seconds_ls leds_seconds_ls (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_leds_seconds_ls_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_seconds_ls_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_seconds_ls_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_seconds_ls_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_seconds_ls_s1_readdata),   //                    .readdata
		.out_port   (leds_seconds_ls_external_connection_export)       // external_connection.export
	);

	cpu_leds_seconds_ls leds_seconds_ms (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_leds_seconds_ms_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_seconds_ms_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_seconds_ms_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_seconds_ms_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_seconds_ms_s1_readdata),   //                    .readdata
		.out_port   (leds_seconds_ms_external_connection_export)       // external_connection.export
	);

	cpu_memoria memoria (
		.clk        (clk_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_memoria_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memoria_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memoria_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memoria_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memoria_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memoria_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memoria_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),      //       .reset_req
		.freeze     (1'b0)                                     // (terminated)
	);

	cpu_pio_key_0 pio_key_0 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_pio_key_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_key_0_s1_readdata), //                    .readdata
		.in_port  (pio_key_0_external_connection_export)     // external_connection.export
	);

	cpu_pio_key_0 pio_key_1 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_pio_key_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_key_1_s1_readdata), //                    .readdata
		.in_port  (pio_key_1_external_connection_export)     // external_connection.export
	);

	cpu_pio_key_0 pio_key_2 (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_pio_key_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_key_2_s1_readdata), //                    .readdata
		.in_port  (pio_key_2_external_connection_export)     // external_connection.export
	);

	cpu_pio_key_3 pio_key_3 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_pio_key_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_key_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_key_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_key_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_key_3_s1_readdata),   //                    .readdata
		.in_port    (pio_key_3_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                   //                 irq.irq
	);

	cpu_pio_switches pio_switches (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_pio_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_switches_s1_readdata), //                    .readdata
		.in_port  (pio_switches_external_connection_export)     // external_connection.export
	);

	cpu_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	cpu_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                             (clk_clk),                                                     //                       clk_0_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                              // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                   (cpu_data_master_address),                                     //                 cpu_data_master.address
		.cpu_data_master_waitrequest               (cpu_data_master_waitrequest),                                 //                                .waitrequest
		.cpu_data_master_byteenable                (cpu_data_master_byteenable),                                  //                                .byteenable
		.cpu_data_master_read                      (cpu_data_master_read),                                        //                                .read
		.cpu_data_master_readdata                  (cpu_data_master_readdata),                                    //                                .readdata
		.cpu_data_master_write                     (cpu_data_master_write),                                       //                                .write
		.cpu_data_master_writedata                 (cpu_data_master_writedata),                                   //                                .writedata
		.cpu_data_master_debugaccess               (cpu_data_master_debugaccess),                                 //                                .debugaccess
		.cpu_instruction_master_address            (cpu_instruction_master_address),                              //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest        (cpu_instruction_master_waitrequest),                          //                                .waitrequest
		.cpu_instruction_master_read               (cpu_instruction_master_read),                                 //                                .read
		.cpu_instruction_master_readdata           (cpu_instruction_master_readdata),                             //                                .readdata
		.cpu_debug_mem_slave_address               (mm_interconnect_0_cpu_debug_mem_slave_address),               //             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                 (mm_interconnect_0_cpu_debug_mem_slave_write),                 //                                .write
		.cpu_debug_mem_slave_read                  (mm_interconnect_0_cpu_debug_mem_slave_read),                  //                                .read
		.cpu_debug_mem_slave_readdata              (mm_interconnect_0_cpu_debug_mem_slave_readdata),              //                                .readdata
		.cpu_debug_mem_slave_writedata             (mm_interconnect_0_cpu_debug_mem_slave_writedata),             //                                .writedata
		.cpu_debug_mem_slave_byteenable            (mm_interconnect_0_cpu_debug_mem_slave_byteenable),            //                                .byteenable
		.cpu_debug_mem_slave_waitrequest           (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),           //                                .waitrequest
		.cpu_debug_mem_slave_debugaccess           (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),           //                                .debugaccess
		.jtag_uart_0_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //   jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                .write
		.jtag_uart_0_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                .read
		.jtag_uart_0_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                .chipselect
		.leds_minutes_ls_s1_address                (mm_interconnect_0_leds_minutes_ls_s1_address),                //              leds_minutes_ls_s1.address
		.leds_minutes_ls_s1_write                  (mm_interconnect_0_leds_minutes_ls_s1_write),                  //                                .write
		.leds_minutes_ls_s1_readdata               (mm_interconnect_0_leds_minutes_ls_s1_readdata),               //                                .readdata
		.leds_minutes_ls_s1_writedata              (mm_interconnect_0_leds_minutes_ls_s1_writedata),              //                                .writedata
		.leds_minutes_ls_s1_chipselect             (mm_interconnect_0_leds_minutes_ls_s1_chipselect),             //                                .chipselect
		.leds_minutes_ms_s1_address                (mm_interconnect_0_leds_minutes_ms_s1_address),                //              leds_minutes_ms_s1.address
		.leds_minutes_ms_s1_write                  (mm_interconnect_0_leds_minutes_ms_s1_write),                  //                                .write
		.leds_minutes_ms_s1_readdata               (mm_interconnect_0_leds_minutes_ms_s1_readdata),               //                                .readdata
		.leds_minutes_ms_s1_writedata              (mm_interconnect_0_leds_minutes_ms_s1_writedata),              //                                .writedata
		.leds_minutes_ms_s1_chipselect             (mm_interconnect_0_leds_minutes_ms_s1_chipselect),             //                                .chipselect
		.leds_seconds_ls_s1_address                (mm_interconnect_0_leds_seconds_ls_s1_address),                //              leds_seconds_ls_s1.address
		.leds_seconds_ls_s1_write                  (mm_interconnect_0_leds_seconds_ls_s1_write),                  //                                .write
		.leds_seconds_ls_s1_readdata               (mm_interconnect_0_leds_seconds_ls_s1_readdata),               //                                .readdata
		.leds_seconds_ls_s1_writedata              (mm_interconnect_0_leds_seconds_ls_s1_writedata),              //                                .writedata
		.leds_seconds_ls_s1_chipselect             (mm_interconnect_0_leds_seconds_ls_s1_chipselect),             //                                .chipselect
		.leds_seconds_ms_s1_address                (mm_interconnect_0_leds_seconds_ms_s1_address),                //              leds_seconds_ms_s1.address
		.leds_seconds_ms_s1_write                  (mm_interconnect_0_leds_seconds_ms_s1_write),                  //                                .write
		.leds_seconds_ms_s1_readdata               (mm_interconnect_0_leds_seconds_ms_s1_readdata),               //                                .readdata
		.leds_seconds_ms_s1_writedata              (mm_interconnect_0_leds_seconds_ms_s1_writedata),              //                                .writedata
		.leds_seconds_ms_s1_chipselect             (mm_interconnect_0_leds_seconds_ms_s1_chipselect),             //                                .chipselect
		.memoria_s1_address                        (mm_interconnect_0_memoria_s1_address),                        //                      memoria_s1.address
		.memoria_s1_write                          (mm_interconnect_0_memoria_s1_write),                          //                                .write
		.memoria_s1_readdata                       (mm_interconnect_0_memoria_s1_readdata),                       //                                .readdata
		.memoria_s1_writedata                      (mm_interconnect_0_memoria_s1_writedata),                      //                                .writedata
		.memoria_s1_byteenable                     (mm_interconnect_0_memoria_s1_byteenable),                     //                                .byteenable
		.memoria_s1_chipselect                     (mm_interconnect_0_memoria_s1_chipselect),                     //                                .chipselect
		.memoria_s1_clken                          (mm_interconnect_0_memoria_s1_clken),                          //                                .clken
		.pio_key_0_s1_address                      (mm_interconnect_0_pio_key_0_s1_address),                      //                    pio_key_0_s1.address
		.pio_key_0_s1_readdata                     (mm_interconnect_0_pio_key_0_s1_readdata),                     //                                .readdata
		.pio_key_1_s1_address                      (mm_interconnect_0_pio_key_1_s1_address),                      //                    pio_key_1_s1.address
		.pio_key_1_s1_readdata                     (mm_interconnect_0_pio_key_1_s1_readdata),                     //                                .readdata
		.pio_key_2_s1_address                      (mm_interconnect_0_pio_key_2_s1_address),                      //                    pio_key_2_s1.address
		.pio_key_2_s1_readdata                     (mm_interconnect_0_pio_key_2_s1_readdata),                     //                                .readdata
		.pio_key_3_s1_address                      (mm_interconnect_0_pio_key_3_s1_address),                      //                    pio_key_3_s1.address
		.pio_key_3_s1_write                        (mm_interconnect_0_pio_key_3_s1_write),                        //                                .write
		.pio_key_3_s1_readdata                     (mm_interconnect_0_pio_key_3_s1_readdata),                     //                                .readdata
		.pio_key_3_s1_writedata                    (mm_interconnect_0_pio_key_3_s1_writedata),                    //                                .writedata
		.pio_key_3_s1_chipselect                   (mm_interconnect_0_pio_key_3_s1_chipselect),                   //                                .chipselect
		.pio_switches_s1_address                   (mm_interconnect_0_pio_switches_s1_address),                   //                 pio_switches_s1.address
		.pio_switches_s1_readdata                  (mm_interconnect_0_pio_switches_s1_readdata),                  //                                .readdata
		.timer_s1_address                          (mm_interconnect_0_timer_s1_address),                          //                        timer_s1.address
		.timer_s1_write                            (mm_interconnect_0_timer_s1_write),                            //                                .write
		.timer_s1_readdata                         (mm_interconnect_0_timer_s1_readdata),                         //                                .readdata
		.timer_s1_writedata                        (mm_interconnect_0_timer_s1_writedata),                        //                                .writedata
		.timer_s1_chipselect                       (mm_interconnect_0_timer_s1_chipselect)                        //                                .chipselect
	);

	cpu_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
